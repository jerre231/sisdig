LIBRARY IEEE;  																				
USE IEEE.STD_LOGIC_1164.ALL;  															
USE IEEE.NUMERIC_STD.ALL;  																

ENTITY LEITOR_TECLA IS
	PORT (
			CLK, RESET: IN  STD_LOGIC;  					-- ENTRADAS DE CLOCK E RESET
			PS2D, PS2C: IN  STD_LOGIC;  					-- ENTRADAS DE DADOS E CLOCK PS2
			LEDS : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);  		-- SAIDA PARA OS LEDS
			TECLOU : OUT STD_LOGIC);  						-- SAIDA PARA INDICAR TECLA PRESSIONADA
END LEITOR_TECLA;

ARCHITECTURE BEHAVIORAL OF LEITOR_TECLA IS

	COMPONENT KB_CODE PORT (
				CLK, RESET: IN  STD_LOGIC;  					-- ENTRADAS DE CLOCK E RESET
				PS2D, PS2C: IN  STD_LOGIC;  					-- ENTRADAS DE DADOS E CLOCK PS2
				RD_KEY_CODE: IN STD_LOGIC;  					-- ENTRADA PARA LER CODIGO DA TECLA
				KEY_CODE: OUT STD_LOGIC_VECTOR(7 DOWNTO 0);     -- SAIDA DO CODIGO DA TECLA
				KB_BUF_EMPTY: OUT STD_LOGIC);  					-- SAIDA INDICANDO BUFFER DO TECLADO VAZIO
			
	END COMPONENT KB_CODE;
	
	TYPE ESTADOS IS (
				EINICIAL,  	-- ESTADO INICIAL
				EMEIO,  	-- ESTADO INTERMEDIARIO
				EFINAL);  	-- ESTADO FINAL
	
	SIGNAL EATUAL : ESTADOS := EINICIAL; 							-- SINAL PARA O ESTADO ATUAL
	SIGNAL EPROXIMO : ESTADOS;  									-- SINAL PARA O PROXIMO ESTADO
	SIGNAL LIBERABUF : STD_LOGIC := '0';  							-- SINAL PARA LIBERAR BUFFER
	SIGNAL KEYREAD : STD_LOGIC_VECTOR (7 DOWNTO 0):= "00000000";  	-- SINAL PARA LEITURA DA TECLA
	SIGNAL KEYBUFFER : STD_LOGIC_VECTOR (7 DOWNTO 0);  				-- SINAL PARA BUFFER DA TECLA
	SIGNAL BUFEMPTY : STD_LOGIC ;  									-- SINAL INDICANDO BUFFER VAZIO
	SIGNAL CLKREDUZIDO : STD_LOGIC := '0';  						-- SINAL DO CLOCK REDUZIDO
	
BEGIN
	KBC: KB_CODE PORT MAP (CLK, RESET, PS2D, PS2C, LIBERABUF, KEYBUFFER, BUFEMPTY);  -- MAPEAMENTO DO COMPONENTE KB_CODE
	LEDS <= KEYREAD;  -- LEDS EXIBEM A TECLA LIDA

	-------------------------------------
	----------REDUTOR DE CLOCK-----------
	-------------------------------------
	PROCESS(CLK)
		VARIABLE CONTAGEM : UNSIGNED (5 DOWNTO 0) := "000000";  	-- VARIAVEL PARA CONTAGEM
		BEGIN
			IF (CLK = '1' AND CLK'EVENT) THEN  						-- SE HOUVER EVENTO DE CLOCK
				IF (CONTAGEM >= 9) THEN  							-- SE A CONTAGEM ATINGIR 9
					CONTAGEM := "000000";  							-- RESETA A CONTAGEM
					CLKREDUZIDO<= NOT CLKREDUZIDO;  				-- INVERTE O CLOCK REDUZIDO
				ELSE
					CONTAGEM := CONTAGEM + 1;  						-- INCREMENTA A CONTAGEM
				END IF;
			END IF;
	END PROCESS;
	
	-------------------------------------
	--------CONTROLE DOS ESTADOS---------
	-------------------------------------
	PROCESS(CLKREDUZIDO, EATUAL, BUFEMPTY)
	BEGIN
		IF (CLKREDUZIDO = '1' AND CLKREDUZIDO'EVENT) THEN  -- SE HOUVER EVENTO DE CLOCK REDUZIDO
			IF EATUAL = EINICIAL THEN  					   -- SE ESTIVER NO ESTADO INICIAL
				IF BUFEMPTY = '0' THEN  				   -- SE O BUFFER NAO ESTIVER VAZIO
					EATUAL <= EMEIO;  					   -- VAI PARA O ESTADO INTERMEDIARIO
				END IF;
			END IF;
			IF EATUAL = EMEIO THEN  					   -- SE ESTIVER NO ESTADO INTERMEDIARIO
				EATUAL <= EFINAL;  						   -- VAI PARA O ESTADO FINAL
			END IF;
			IF EATUAL = EFINAL THEN  					   -- SE ESTIVER NO ESTADO FINAL
				EATUAL <= EINICIAL;  					   -- VOLTA PARA O ESTADO INICIAL
			END IF;
		END IF;
	END PROCESS;
	
	-- PROCESSO PARA A��ES EM CADA ESTADO
	PROCESS(CLKREDUZIDO)
	BEGIN
		IF EATUAL = EINICIAL THEN  		-- SE ESTIVER NO ESTADO INICIAL
			LIBERABUF <= '0';  			-- NAO LIBERA O BUFFER
		END IF;
		IF EATUAL = EMEIO THEN  		-- SE ESTIVER NO ESTADO INTERMEDIARIO
			KEYREAD <= KEYBUFFER;  		-- LE O BUFFER DA TECLA
		END IF;
		IF EATUAL = EFINAL THEN  		-- SE ESTIVER NO ESTADO FINAL
			LIBERABUF <= '1';  			-- LIBERA O BUFFER
		END IF;
	END PROCESS;
END BEHAVIORAL;

